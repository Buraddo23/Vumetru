library verilog;
use verilog.vl_types.all;
entity top_tb is
    generic(
        delay           : integer := 128
    );
end top_tb;
