library verilog;
use verilog.vl_types.all;
entity clk_gen_tb is
end clk_gen_tb;
