library verilog;
use verilog.vl_types.all;
entity img_tb is
end img_tb;
