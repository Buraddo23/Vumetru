library verilog;
use verilog.vl_types.all;
entity uart_tb is
    generic(
        delay           : integer := 32
    );
end uart_tb;
