library verilog;
use verilog.vl_types.all;
entity top_clk_gen_tb is
end top_clk_gen_tb;
